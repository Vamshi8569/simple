import uvm_pkg::*;
`include "uvm_macros.svh"

`include "mem_tx.sv"
`include "mem_seq.sv"
`include "mem_sqr.sv"
`include "mem_driver.sv"
`include "mem_agent.sv"
`include "mem_env.sv"
`include "mem_test.sv"
`include "top.sv"

